package v10_filter_parameters;

	parameter k_var10=4'd10;
	parameter l_var10=3'd6;
	parameter M_var10=5'd16;
	parameter M_length_var10=3'd4;
	
endpackage
