package v10_filter_parameters;

	parameter k_var10=4'd10;
	parameter l_var10=3'd6;
	parameter M_var10=4'd15;
	parameter Mw_var10=3'd4;
	
endpackage
