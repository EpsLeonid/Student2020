package registr_parameter;
parameter width=8;
endpackage
