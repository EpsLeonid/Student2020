package v9_parameter;
	parameter l_9 = 6;
	parameter k_9 = 13;
	parameter m1 = 15;
	parameter m2 = 1;
endpackage