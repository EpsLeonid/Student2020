package Register_param;
	parameter  bus_width=4'd8;
endpackage