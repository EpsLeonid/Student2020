package reg_param;

	localparam bus_width=4'd8;
	
endpackage