module qqq(A,B,C);
				
input A;
input B;
output C;
assign C=A*B;
endmodule 