package v8_param;

	parameter k_var8=3'd7;
	parameter l_var8=3'd7;
	parameter M_var8=5'd16;
	
endpackage