package v9_parameters;

parameter v9_k=13;
parameter v9_l=6;
parameter v9_m1=15;
parameter v9_m2=1;
parameter SIZE = 20;

endpackage
