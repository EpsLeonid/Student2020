package v10_filter_parameters;

parameter k_10=10;
parameter l_10=6;
parameter M_10=16;
endpackage