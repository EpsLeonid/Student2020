package v5_param;

	parameter k_var5=3'd6;
	parameter l_var5=3'd6;
	parameter M_var5=7'd16;
	parameter M_dig_var5=3'd4;
	
endpackage
