package registr_parameter;
parameter size=8;
endpackage 