package v10_filter_parameters;

	parameter k_var7=4'd10;
	parameter l_var7=3'd6;
	parameter M_var7=5'd16;
	parameter M_length_var7=3'd4;
	
endpackage
