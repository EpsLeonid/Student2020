module multiply(output C,
				input A,B
				);
				
	and AND1(C, A,B);

endmodule