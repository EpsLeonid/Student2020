module ABC(input [3:0]B, C,
				output [7:0]A);
	assign A = B * C;
	
	endmodule
				