package v4_filter_parameters;
parameter K=9;
parameter L=5;
parameter M=16;
endpackage