package v10_filter_parameters;

	parameter   k_v10=4'd10, 
				l_v10=3'd6,
				M_v10=5'd16,
				M_length_v10=3'd4;	
endpackage
