package register_parameter;
parameter size=8;
endpackage