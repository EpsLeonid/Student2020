package v3_filter_parameters;


parameter v3_k=11;
parameter v3_l=5;
parameter v3_m1=16;
parameter v3_m2=1;
parameter SIZE = 20;
endpackage
