package v7_param;

	parameter k_var7=4'd10;
	parameter l_var7=3'd5;
	parameter M_var7=4'd15;
	parameter M_length_var7=3'd4;
	
endpackage