package Parametrs_reg;
parameter input_size=8;
parameter output_size=16;
endpackage
