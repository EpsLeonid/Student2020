package task3_parameter;
parameter size=8;
endpackage