package ABC_parameter;
parameter lenght=8;
endpackage