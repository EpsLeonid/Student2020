package parameters_v2;
	parameter M = 16;
	parameter k = 5;
	parameter l = 5;
endpackage