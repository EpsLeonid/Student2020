package Bits;

	parameter SIZE = 8;

	
endpackage
