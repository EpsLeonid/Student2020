package v1_param;

	parameter k_var1=4'd8;
	parameter l_var1=3'd5;
	parameter M_var1=5'd16;
	
endpackage