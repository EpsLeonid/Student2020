package v3_filter_parameters;

parameter m1=16;
parameter m2=1;
parameter k=11;
parameter l=5;
parameter SIZE_ADC_DATA = 20;

endpackage
