package v5_param;

parameter M_5 = 16;
parameter l_5 = 6;
parameter k_5 = 6;
endpackage