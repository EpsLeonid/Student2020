module zadanie1(A,B,C);

input wire A;
input wire B;
output C;

assign C=A*B;

endmodule
