package v5_param;

parameter k=16;
parameter l=6;
parameter m=6;
endpackage