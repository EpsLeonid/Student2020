package parameter1;
parameter width=8;
parameter a=width*width;
parameter b=a+width;
endpackage
