module task1(A,B,C);
input wire A, B;
output reg C=1'b0;

assign C=A*B;

endmodule