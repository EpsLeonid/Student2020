package v6_parameters;

parameter v6_k=13;
parameter v6_l=6;
parameter v6_m1=16;
parameter v6_m2=1;


endpackage
