package Bits;

	parameter SIZE = 4;

	
endpackage