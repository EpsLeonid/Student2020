package v8_param;

	parameter k_var8=3'd7;
	parameter l_var8=3'd7;
	parameter M_var8=4'd15;
	parameter M_dig_var8=3'd4;
	
endpackage