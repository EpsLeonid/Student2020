package v10_filter_parameters;

	parameter   k_v10=4'd10; 
	parameter	l_v10=3'd6;
	parameter	M_v10=5'd16;
endpackage
